    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   SaveData   clases	variablesobjetosreferenciasconsolauSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   	   	   	   	   	      uSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  
ClaseSav[]   	            xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  VariableSav[]   		              ~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	
                 	
              System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	                   ClaseSav   	   	           VariableSav   
                N<#7D81CF>clase1</color> <#63A7A6>var2</color> = new <#7D81CF>clase1</color>();   N<#7D81CF>clase1</color> <#63A7A6>var2</color> = new <#7D81CF>clase1</color>();   N<#7D81CF>clase1</color> <#1D2F53>var1</color> = new <#7D81CF>clase1</color>();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   ClaseSav   nombrecolor	atributosmetodosxSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]      clase1	   	   	         .0�>�&?��O?   xSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  AtributoSav[]   	            vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  MetodoSav[]   	                   AtributoSav   	             	MetodoSav   	       AtributoSav   nombretipo
proteccion   !   x"   int#   Public    	MetodoSav   nombre   $   Read�'?(o&?&          AtributoSav   	(   '          	MetodoSav   	)   (   AtributoSav   nombretipo
proteccion   *   x+   int,   Public)   	MetodoSav   nombre   -   Read