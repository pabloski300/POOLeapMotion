    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   SaveData   clases	variablesobjetosuSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   	   	   	      uSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  
ClaseSav[]   	            xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  VariableSav[]   	            ~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	                   ClaseSav   		             VariableSav   	
                         	   ClaseSav   nombrecolor	atributosmetodosxSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]      clase	   	   	   
   VariableSav   clasenombrecolor   	      var	         J�_?F�X?��:?   xSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  AtributoSav[]   	              vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  MetodoSav[]   	               ��a?j��>��P?           AtributoSav             	MetodoSav   	      	MetodoSav   nombre      
MetodoRead    AtributoSav              	MetodoSav             AtributoSav   	             	MetodoSav   	      AtributoSav   nombretipo
proteccion      x   int   Public   	MetodoSav   nombre       
MetodoRead