    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   SaveData   clases	variablesobjetosreferenciasconsolauSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   	   	   	   	   	      uSystem.Collections.Generic.List`1[[ClaseSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  
ClaseSav[]   	            xSystem.Collections.Generic.List`1[[VariableSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  VariableSav[]   		            ~System.Collections.Generic.List`1[[System.Int32, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	
               	            System.Collections.Generic.List`1[[System.String, mscorlib, Version=4.0.0.0, Culture=neutral, PublicKeyToken=b77a5c561934e089]]   _items_size_version  	                   ClaseSav   	   	   	          VariableSav   	   	   
                           ����                    var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   var1.Read();   -<#7D81CF>clase1</color> <#17E14E>var</color>;   new <#7D81CF>clase1</color>();   .<#A20236>clase2</color> <#BDA79F>var2</color>;   new <#A20236>clase2</color>();   6<#BDA79F>var2</color> = new <#A20236>clase2</color>();    <#BDA79F>var2</color>.Sub(0, 0);   ClaseSav   nombrecolor	atributosmetodosxSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]      clase1	   	   	          !   clase2	"   	#   	$      VariableSav   clasenombrecolor   	   &   var	'         	!   )   var2	*         .0�>�&?��O?   xSystem.Collections.Generic.List`1[[AtributoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  AtributoSav[]   	+             vSystem.Collections.Generic.List`1[[MetodoSav, Assembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null]]   _items_size_version  MetodoSav[]   	,         "      �"? <`�X>#      	-         $       	.         '      ���=LNb?���>*      \*>?:�'?�
 ?+          AtributoSav   	/   ,          	MetodoSav   	0   -          AtributoSav   	1   .          	MetodoSav   	2   /   AtributoSav   nombretipo
proteccion   3   x4   int5   Public0   	MetodoSav   nombre   6   Read1   /   7   x8   bool	5   2   0   :   Sub